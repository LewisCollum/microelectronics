.subckt inverter vDD input output
.param sourceLength=1u sourceWidth=16u sinkLength=1u sinkWidth=8u

mSource output input vDD sourceBody source
+ L = sourceLength
+ W = sourceWidth

mSink output input 0 sinkBody sink
+ L = sinkLength
+ W = sinkWidth
.ends


.model source pmos
+ kp = 0.08m
+ vto = -1
+ lambda = 0.2
+ cbd = 100fF
+ cbs = 100fF
+ tox = 50nm 

.model sink nmos
+ kp = 0.18m
+ vto = 1
+ lambda = 0.2
+ cbd = 100fF
+ cbs = 100fF
+ tox = 50nm
